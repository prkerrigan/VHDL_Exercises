ENTITY test_bench4 IS
END ENTITY test_bench4;


